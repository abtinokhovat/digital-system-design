library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity generator is
 port();
end generator;
 
architecture behavior of generator is
begin
end behavior;

