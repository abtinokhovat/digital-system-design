library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity checker is
 port();
end checker;
 
architecture behavior of checker is
begin
end behavior;

